--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   12:58:08 10/29/2018
-- Design Name:   
-- Module Name:   C:/Users/Alejandro ramirez/Desktop/xilink/FFR/tb_FFR.vhd
-- Project Name:  FFR
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: FFR
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_FFR IS
END tb_FFR;
 
ARCHITECTURE behavior OF tb_FFR IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT FFR
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         d : IN  std_logic_vector(1 downto 0);
         q : OUT  std_logic_vector(1 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';
   signal d : std_logic_vector(1 downto 0) := (others => '0');

 	--Outputs
   signal q : std_logic_vector(1 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: FFR PORT MAP (
          clk => clk,
          rst => rst,
          d => d,
          q => q
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		

      -- hold reset state for 100 ns.
      wait for 100 ns;	
		
		wait for 4 ns;
		d <= "10";
		wait for 4 ns;
		d <= "11";
		wait for 15 ns;
		d <= "10";
		wait for 1 ns;
		d <= "11";
		wait for 15 ns;
		rst <= '1';

      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
